ELF          *            �
     4     (  	             �/�/ �/�/�/�/C��/C�"O� �dH$�A�@	 �.@��dH$�=�B	 �-=��dH$�9�C	 �,:۲dH$�5�E	 �+�h6�7ن�g6�y�fg�dH4�H	 �dH.2�H-�dH,+�c8#��b("��a!� �6 �)&O�n�m�l�k�j�i �h	 	 	 	 � �ܢ)�dH$��K	 �,۲dH$��M	 �+ْdH$��N	 �)؂dH$�	�@	 �(�e��
�V�c9�b'�lů�                          �       �  0�  	 	 	 	 	 	 	 	 	 	 	 	 �/ �/wئ/wж/"O" H	  ���&O�k�j�i �hp� �p�$֕�o�	�	�	�	�	��2g��/�ZH �-�,��,����ZF-�v���b�ZFr�B�vG6*�w��w-�:�wZ��w��sirj\9�)b�qSr�1B�rR"s[�sk{w*��i��\9w:�wZ��wtZ�) w�S1�R"�ZǏ�x8��ZHN� �N� 炙 � � ��s`Bc-@�(Rb32��cbRc�2&Rc32br!Rc32b r"Ba�1���!�wr!=wBbs`�wh&@2qBa�w�1����wrwR`�scBbC<0<2pr��R`<0QR`<0b!r%R`<0QBb<2�76`�scs4�BasbB-�28E�r>wq�wBasb�vB2v3g�76���x.�g8�� {�G��Bh|8�I��I	 � �%�&O `b                 �A  �<   =���<  �A��*<             T   ���	 	 	 	 	 	 	 	 	 	 	 	 	 	 ���s	 	 	 	 	 	 	 	 	 	 	 	 	 q�R`	 	 	 	 	 	 	 	 	 	 	 	 	 	 P�Bb	 	 	 	 	 	 	 	 	 	 	 	 	 	 �/�//�/�/�/�/�/��q��"Oq�חabc7sShx�`� ��C0��0�x�Sh
�"`p"x��x*�"jz�"x�H:�"k{��"x��x�(z�"dtB"x�j�"n~�"x�Z�"m}�"x�J�"l|��"FȏShR���R�镕bdQ�Q�HL5L� 排 �Rc����,3��3aL�	�<7�D��c`�@0�B�B)�ZBZBx�\6-�c`B�qsc�@��0s�0�^���B��q��B)ZB8�\6-�c`B�qsc�@��0 s��0�^���B��q��B)ZB8�\6-�c`B�$qsc�@��00sl�0�^���B`��qZB8�4q-��xB�@w�(\6����0�^�z�q� ��>�����d�x�f�4�e�6�4K�6�g�dw�f y�e|4|6�4K�6�(�&O���n�m�l�k�j�i �h� ^�4 @	 RI7               @�  ��>��Y?       	 	 	 	 	 	 	 	 	 	 	 	 	 	 ��B)	 	 	 	 	 	 	 	 	 	 	 	 	 	 {�ZB	 	 	 	 	 	 	 	 	 	 	 	 	 	 U�ZB	 	 	 	 	 	 	 	 	 	 	 	 	 	 �/�/�/ �/��/"Oܒ � �dH$��@	 �,۲dH$��B	 �+ڢdH$��C	 �*؂dH$��E	 �(�`��i��gw�fh&O�l�k�j�i �h                         	 	 	 	 	 	 	 	 � ��"O�2%�2$2"2 �2 &O  �	                  	 	 	 	 	 	 �/�/�/ �/��/"Oܒ � �dH$��@	 �,۲dH$��B	 �+ڢdH$��C	 �*؂dH$��E	 �(�`��i ���gw�fh&O�l�k�j�i �h	                          	 	 	 	 	 	 �Ce"O"` ���C	 �@	  �&O 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 ���        T      	 	 	 	 	 	 "O&O  �	 	 	 	 	 	 	 	 	 	 	 	 �"O"` � ��	�����@�� �&O 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 ���      �Bfff?        T   	 	 "O&O c`	 	 	 	 	 	 	 	 	 	 	 	 "O�&O 	 	 (   	 	 	 	 	 	 	 	 fft-vlr FFT-VLR Vincent Penne Benjamin Gerard   Virtual Landscape Reality based on Fast Fourier Transform              b     b                      VIS          0          `  �  `  �     `  �   GCC: (GNU) 3.0.4 �ޭ� .symtab .strtab .shstrtab .rela.text .rodata .rela.data .bss .comment .stack                                                       @    	                                �  d  
            &             `	  l                  3             �	  d                  .              H  �   
            9             0
  �                  >              0
                    G             B
                                  F
  N                                t                	              �  ]                                                                                                                                                            ��              #              0              8    	       A              M              T               _free _MtxCopy _ready _FaceNormal _MtxIdentity _malloc _ko_main _DrawObject _fft_F _memmove      	               $        (        ,        0        4        <        D        H  	      L        P        l        p        t        x        |        �        �        �        �        �           
      �  	      �        �                                         @  	      D        H        L        P        �  	      �        �        �        �        �        �        D  	      H        L        P        �  	      �        �        �        	                  4         8         <         D         H         L         P         T         X         \         `         